module registerFile
(
	input [4:0] rs1,
	input [4:0] rs2,
	input [4:0] rd,
	input [63:0] Write_Data,
	input clk, reset, Reg_Write,
	output reg [63:0] Read_Data1,
	output reg [63:0] Read_Data2
	
);

reg [63:0] register [17:0] ;
	initial
	begin
	register[0] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000;
	register[1] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001;
	register[2] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0010;
	register[3] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0011;
	register[4] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0100;
	register[5] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0101;
	register[6] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0110;
	register[7] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0111;
	register[8] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1000;
	register[9] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1001;
	register[10] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1010;
	register[11] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1011;
	register[12] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1100;
	register[13] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1101;
	register[14] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1110;
	register[15] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_1111;
	register[16] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0000;
	register[17] = 64'b 0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0000_0001_0001;
	end

	always@(posedge clk or posedge reset )
		begin
		Read_Data1 = register[rs1];
		Read_Data2 = register[rs2];
			if (Reg_Write == 1)
				register[rd] = Write_Data;
				
			if(reset)
				begin
				Read_Data1 = 64'd0;
				Read_Data2 = 64'd0;
				end
		end
endmodule 